//----------------------------------//
// Breakout Files
// score.v
// David J. Morvay
// ECEN 4856
// Fall 2020
//----------------------------------//

module score(clk, reset, score, pix_x, pix_y, ball_x_r, ball_x_l, ball_y_t, ball_y_b, moveD, moveL, moveR, score_ON_R, score_ON_RM, score_ON_LM, score_ON_L);
input clk, reset;
input [15:0] score;
input [10:0] pix_x, pix_y, ball_x_r, ball_x_l, ball_y_t, ball_y_b;
output moveD, moveL, moveR, score_ON_R, score_ON_RM, score_ON_LM, score_ON_L;


localparam NUM_SIZE = 32;
//-------------------------------------------------------------------------------------------------------------//
// Right Number

// number left, right boundary
wire [10:0] NUM_x_l_1 = 432;
wire [10:0] NUM_x_r_1 = NUM_x_l_1 + NUM_SIZE - 1;
// number top, bottom boundary 
wire [10:0] NUM_y_t_1 = 565; 
wire [10:0] NUM_y_b_1 = NUM_y_t_1 + NUM_SIZE - 1;
reg rom_bit_1;

//------------------------------------//
// Number 0
wire [4:0] rom_addr0_1, rom_col0_1;
reg [31:0] rom_data0_1;

// number image ROM
always @*
case (rom_addr0_1)
	5'h0: rom_data0_1 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data0_1 =   32'b10000000_00000000_00000000_00000000;	//   *                              *
	5'h2: rom_data0_1 =   32'b10000000_00000000_00000000_00000000;	//   *                              *
	5'h3: rom_data0_1 =   32'b10000000_00011111_11111000_00000000;	//   *          **********          *
	5'h4: rom_data0_1 =   32'b10000000_00111111_11111100_00000000;	//   *         ************         *
	5'h5: rom_data0_1 =   32'b10000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h6: rom_data0_1 =   32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h7: rom_data0_1 =   32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h8: rom_data0_1 =   32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h9: rom_data0_1 =   32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hA: rom_data0_1 =   32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hB: rom_data0_1 =   32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hC: rom_data0_1 =   32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hD: rom_data0_1 =   32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hE: rom_data0_1 =   32'b10000000_01000000_00000010_00000000;	//   *        *            *        *
	5'hF: rom_data0_1 =   32'b10000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h10: rom_data0_1 =  32'b10000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h11: rom_data0_1 =  32'b10000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h12: rom_data0_1 =  32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h13: rom_data0_1 =  32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h14: rom_data0_1 =  32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h15: rom_data0_1 =  32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h16: rom_data0_1 =  32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h17: rom_data0_1 =  32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h18: rom_data0_1 =  32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h19: rom_data0_1 =  32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h1A: rom_data0_1 =  32'b10000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h1B: rom_data0_1 =  32'b10000000_00111111_11111100_00000000;	//   *         ************         *
	5'h1C: rom_data0_1 =  32'b10000000_00011111_11111000_00000000;	//   *          **********          *
	5'h1D: rom_data0_1 =  32'b10000000_00000000_00000000_00000000; 	//   *				    *
	5'h1E: rom_data0_1 =  32'b10000000_00000000_00000000_00000000; 	//   *				    *
	5'h1F: rom_data0_1 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr0_1 = pix_y[4:0] - NUM_y_t_1[4:0];
assign rom_col0_1 = pix_x[4:0] - NUM_x_l_1[4:0];

//------------------------------------//
// Number 1
wire [4:0] rom_addr1_1, rom_col1_1;
reg [31:0] rom_data1_1;

// number image ROM
always @*
case (rom_addr1_1)
	5'h0: rom_data1_1 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data1_1 =   32'b10000000_00000000_00000000_00000000;	//   *                              *
	5'h2: rom_data1_1 =   32'b10000000_00000000_00000000_00000000;	//   *                              *
	5'h3: rom_data1_1 =   32'b10000000_00000000_00000000_00000000;	//   *                              *
	5'h4: rom_data1_1 =   32'b10000000_00000000_00000000_00000000;	//   *                              *
	5'h5: rom_data1_1 =   32'b10000000_01000000_00000000_00000000;	//   *        *                     *
	5'h6: rom_data1_1 =   32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h7: rom_data1_1 =   32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h8: rom_data1_1 =   32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h9: rom_data1_1 =   32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'hA: rom_data1_1 =   32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'hB: rom_data1_1 =   32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'hC: rom_data1_1 =   32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'hD: rom_data1_1 =   32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'hE: rom_data1_1 =   32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'hF: rom_data1_1 =   32'b10000000_01000000_00000000_00000000;	//   *        *                     *
	5'h10: rom_data1_1 =  32'b10000000_01000000_00000000_00000000;	//   *        *                     *
	5'h11: rom_data1_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h12: rom_data1_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h13: rom_data1_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h14: rom_data1_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h15: rom_data1_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h16: rom_data1_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h17: rom_data1_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h18: rom_data1_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h19: rom_data1_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h1A: rom_data1_1 =  32'b10000000_01000000_00000000_00000000;	//   *        *                     *
	5'h1B: rom_data1_1 =  32'b10000000_00000000_00000000_00000000;	//   *                              *
	5'h1C: rom_data1_1 =  32'b10000000_00000000_00000000_00000000;	//   *                              *
	5'h1D: rom_data1_1 =  32'b10000000_00000000_00000000_00000000; 	//   *				    *
	5'h1E: rom_data1_1 =  32'b10000000_00000000_00000000_00000000; 	//   *				    *
	5'h1F: rom_data1_1 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr1_1 = pix_y[4:0] - NUM_y_t_1[4:0];
assign rom_col1_1 = pix_x[4:0] - NUM_x_l_1[4:0];

//------------------------------------//
// Number 2
wire [4:0] rom_addr2_1, rom_col2_1;
reg [31:0] rom_data2_1;

// number image ROM
always @*
case (rom_addr2_1)
	5'h0: rom_data2_1 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data2_1 =   32'b10000000_00000000_00000000_00000000;	//   *                              *
	5'h2: rom_data2_1 =   32'b10000000_00000000_00000000_00000000;	//   *                              *
	5'h3: rom_data2_1 =   32'b10000000_00011111_11111000_00000000;	//   *          **********          *
	5'h4: rom_data2_1 =   32'b10000000_00111111_11111100_00000000;	//   *         ************         *
	5'h5: rom_data2_1 =   32'b10000000_01000000_00000000_00000000;	//   *        *                     *
	5'h6: rom_data2_1 =   32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h7: rom_data2_1 =   32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h8: rom_data2_1 =   32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h9: rom_data2_1 =   32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'hA: rom_data2_1 =   32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'hB: rom_data2_1 =   32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'hC: rom_data2_1 =   32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'hD: rom_data2_1 =   32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'hE: rom_data2_1 =   32'b10000000_01000000_00000000_00000000;	//   *        *                     *
	5'hF: rom_data2_1 =   32'b10000000_00111111_11111100_00000000;	//   *         ************         *
	5'h10: rom_data2_1 =  32'b10000000_00111111_11111100_00000000; 	//   *         ************         *
	5'h11: rom_data2_1 =  32'b10000000_00000000_00000010_00000000;	//   *                     *        *
	5'h12: rom_data2_1 =  32'b10000000_00000000_00000011_00000000;	//   *                     **       *
	5'h13: rom_data2_1 =  32'b10000000_00000000_00000011_00000000;	//   *                     **       *
	5'h14: rom_data2_1 =  32'b10000000_00000000_00000011_00000000;	//   *                     **       *
	5'h15: rom_data2_1 =  32'b10000000_00000000_00000011_00000000;	//   *                     **       *
	5'h16: rom_data2_1 =  32'b10000000_00000000_00000011_00000000;	//   *                     **       *
	5'h17: rom_data2_1 =  32'b10000000_00000000_00000011_00000000;	//   *                     **       *
	5'h18: rom_data2_1 =  32'b10000000_00000000_00000011_00000000;	//   *                     **       *
	5'h19: rom_data2_1 =  32'b10000000_00000000_00000011_00000000;	//   *                     **       *
	5'h1A: rom_data2_1 =  32'b10000000_00000000_00000010_00000000;	//   *                     *        *
	5'h1B: rom_data2_1 =  32'b10000000_00111111_11111100_00000000;	//   *         ************         *
	5'h1C: rom_data2_1 =  32'b10000000_00011111_11111000_00000000;	//   *          **********          *
	5'h1D: rom_data2_1 =  32'b10000000_00000000_00000000_00000000; 	//   *				    *
	5'h1E: rom_data2_1 =  32'b10000000_00000000_00000000_00000000; 	//   *				    *
	5'h1F: rom_data2_1 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr2_1 = pix_y[4:0] - NUM_y_t_1[4:0];
assign rom_col2_1 = pix_x[4:0] - NUM_x_l_1[4:0];

//------------------------------------//
// Number 3
wire [4:0] rom_addr3_1, rom_col3_1;
reg [31:0] rom_data3_1;

// number image ROM
always @*
case (rom_addr3_1)
	5'h0: rom_data3_1 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data3_1 =   32'b10000000_00000000_00000000_00000000;	//   *                              *
	5'h2: rom_data3_1 =   32'b10000000_00000000_00000000_00000000;	//   *                              *
	5'h3: rom_data3_1 =   32'b10000000_00011111_11111000_00000000;	//   *          **********          *
	5'h4: rom_data3_1 =   32'b10000000_00111111_11111100_00000000;	//   *         ************         *
	5'h5: rom_data3_1 =   32'b10000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h6: rom_data3_1 =   32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h7: rom_data3_1 =   32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h8: rom_data3_1 =   32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h9: rom_data3_1 =   32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'hA: rom_data3_1 =   32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'hB: rom_data3_1 =   32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'hC: rom_data3_1 =   32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'hD: rom_data3_1 =   32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'hE: rom_data3_1 =   32'b10000000_01000000_00000000_00000000;	//   *        *                     *
	5'hF: rom_data3_1 =   32'b10000000_00111111_11111100_00000000;	//   *         ************         *
	5'h10: rom_data3_1 =  32'b10000000_00111111_11111100_00000000; 	//   *         ************         *
	5'h11: rom_data3_1 =  32'b10000000_01000000_00000000_00000000;	//   *        *                     *
	5'h12: rom_data3_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h13: rom_data3_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h14: rom_data3_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h15: rom_data3_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h16: rom_data3_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h17: rom_data3_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h18: rom_data3_1 =  32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h19: rom_data3_1 =  32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h1A: rom_data3_1 =  32'b10000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h1B: rom_data3_1 =  32'b10000000_00111111_11111100_00000000;	//   *         ************         *
	5'h1C: rom_data3_1 =  32'b10000000_00011111_11111000_00000000;	//   *          **********          *
	5'h1D: rom_data3_1 =  32'b10000000_00000000_00000000_00000000; 	//   *				    *
	5'h1E: rom_data3_1 =  32'b10000000_00000000_00000000_00000000; 	//   *				    *
	5'h1F: rom_data3_1 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr3_1 = pix_y[4:0] - NUM_y_t_1[4:0];
assign rom_col3_1 = pix_x[4:0] - NUM_x_l_1[4:0];

//------------------------------------//
// Number 4
wire [4:0] rom_addr4_1, rom_col4_1;
reg [31:0] rom_data4_1;

// number image ROM
always @*
case (rom_addr4_1)
	5'h0: rom_data4_1 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data4_1 =   32'b10000000_00000000_00000000_00000000;	//   *                              *
	5'h2: rom_data4_1 =   32'b10000000_00000000_00000000_00000000;	//   *                              *
	5'h3: rom_data4_1 =   32'b10000000_00000000_00000000_00000000;	//   *                              *
	5'h4: rom_data4_1 =   32'b10000000_00000000_00000000_00000000;	//   *                              *
	5'h5: rom_data4_1 =   32'b10000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h6: rom_data4_1 =   32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h7: rom_data4_1 =   32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h8: rom_data4_1 =   32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h9: rom_data4_1 =   32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hA: rom_data4_1 =   32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hB: rom_data4_1 =   32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hC: rom_data4_1 =   32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hD: rom_data4_1 =   32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hE: rom_data4_1 =   32'b10000000_01000000_00000010_00000000;	//   *        *            *        *
	5'hF: rom_data4_1 =   32'b10000000_00111111_11111100_00000000;	//   *         ************         *
	5'h10: rom_data4_1 =  32'b10000000_00111111_11111100_00000000; 	//   *         ************         *
	5'h11: rom_data4_1 =  32'b10000000_01000000_00000000_00000000;	//   *        *                     *
	5'h12: rom_data4_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h13: rom_data4_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h14: rom_data4_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h15: rom_data4_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h16: rom_data4_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h17: rom_data4_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h18: rom_data4_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h19: rom_data4_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h1A: rom_data4_1 =  32'b10000000_01000000_00000000_00000000;	//   *        *                     *
	5'h1B: rom_data4_1 =  32'b10000000_00000000_00000000_00000000; 	//   *				    *
	5'h1C: rom_data4_1 =  32'b10000000_00000000_00000000_00000000; 	//   *				    *
	5'h1D: rom_data4_1 =  32'b10000000_00000000_00000000_00000000; 	//   *				    *
	5'h1E: rom_data4_1 =  32'b10000000_00000000_00000000_00000000; 	//   *				    *
	5'h1F: rom_data4_1 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr4_1 = pix_y[4:0] - NUM_y_t_1[4:0];
assign rom_col4_1 = pix_x[4:0] - NUM_x_l_1[4:0];

//------------------------------------//
// Number 5
wire [4:0] rom_addr5_1, rom_col5_1;
reg [31:0] rom_data5_1;

// number image ROM
always @*
case (rom_addr5_1)
	5'h0: rom_data5_1 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data5_1 =   32'b10000000_00000000_00000000_00000000;	//   *                              *
	5'h2: rom_data5_1 =   32'b10000000_00000000_00000000_00000000;	//   *                              *
	5'h3: rom_data5_1 =   32'b10000000_00011111_11111000_00000000;	//   *          **********          *
	5'h4: rom_data5_1 =   32'b10000000_00111111_11111100_00000000;	//   *         ************         *
	5'h5: rom_data5_1 =   32'b10000000_00000000_00000010_00000000;	//   *                     *        *
	5'h6: rom_data5_1 =   32'b10000000_00000000_00000011_00000000;	//   *                     **       *
	5'h7: rom_data5_1 =   32'b10000000_00000000_00000011_00000000;	//   *                     **       *
	5'h8: rom_data5_1 =   32'b10000000_00000000_00000011_00000000;	//   *                     **       *
	5'h9: rom_data5_1 =   32'b10000000_00000000_00000011_00000000;	//   *                     **       *
	5'hA: rom_data5_1 =   32'b10000000_00000000_00000011_00000000;	//   *                     **       *
	5'hB: rom_data5_1 =   32'b10000000_00000000_00000011_00000000;	//   *                     **       *
	5'hC: rom_data5_1 =   32'b10000000_00000000_00000011_00000000;	//   *                     **       *
	5'hD: rom_data5_1 =   32'b10000000_00000000_00000011_00000000;	//   *                     **       *
	5'hE: rom_data5_1 =   32'b10000000_00000000_00000010_00000000;	//   *                     *        *
	5'hF: rom_data5_1 =   32'b10000000_00111111_11111100_00000000;	//   *         ************         *
	5'h10: rom_data5_1 =  32'b10000000_00111111_11111100_00000000; 	//   *         ************         *
	5'h11: rom_data5_1 =  32'b10000000_01000000_00000000_00000000;	//   *        *                     *
	5'h12: rom_data5_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h13: rom_data5_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h14: rom_data5_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h15: rom_data5_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h16: rom_data5_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h17: rom_data5_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h18: rom_data5_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h19: rom_data5_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h1A: rom_data5_1 =  32'b10000000_01000000_00000000_00000000;	//   *        *                     *
	5'h1B: rom_data5_1 =  32'b10000000_00111111_11111100_00000000;	//   *         ************         *
	5'h1C: rom_data5_1 =  32'b10000000_00011111_11111000_00000000;	//   *          **********          *
	5'h1D: rom_data5_1 =  32'b10000000_00000000_00000000_00000000; 	//   *				    *
	5'h1E: rom_data5_1 =  32'b10000000_00000000_00000000_00000000; 	//   *				    *
	5'h1F: rom_data5_1 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr5_1 = pix_y[4:0] - NUM_y_t_1[4:0];
assign rom_col5_1 = pix_x[4:0] - NUM_x_l_1[4:0];

//------------------------------------//
// Number 6
wire [4:0] rom_addr6_1, rom_col6_1;
reg [31:0] rom_data6_1;

// number image ROM
always @*
case (rom_addr6_1)
	5'h0: rom_data6_1 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data6_1 =   32'b10000000_00000000_00000000_00000000;	//   *                              *
	5'h2: rom_data6_1 =   32'b10000000_00000000_00000000_00000000;	//   *                              *
	5'h3: rom_data6_1 =   32'b10000000_00011111_11111000_00000000;	//   *          **********          *
	5'h4: rom_data6_1 =   32'b10000000_00111111_11111100_00000000;	//   *         ************         *
	5'h5: rom_data6_1 =   32'b10000000_00000000_00000010_00000000;	//   *                     *        *
	5'h6: rom_data6_1 =   32'b10000000_00000000_00000011_00000000;	//   *                     **       *
	5'h7: rom_data6_1 =   32'b10000000_00000000_00000011_00000000;	//   *                     **       *
	5'h8: rom_data6_1 =   32'b10000000_00000000_00000011_00000000;	//   *                     **       *
	5'h9: rom_data6_1 =   32'b10000000_00000000_00000011_00000000;	//   *                     **       *
	5'hA: rom_data6_1 =   32'b10000000_00000000_00000011_00000000;	//   *                     **       *
	5'hB: rom_data6_1 =   32'b10000000_00000000_00000011_00000000;	//   *                     **       *
	5'hC: rom_data6_1 =   32'b10000000_00000000_00000011_00000000;	//   *                     **       *
	5'hD: rom_data6_1 =   32'b10000000_00000000_00000011_00000000;	//   *                     **       *
	5'hE: rom_data6_1 =   32'b10000000_00000000_00000010_00000000;	//   *                     *        *
	5'hF: rom_data6_1 =   32'b10000000_00111111_11111100_00000000;	//   *         ************         *
	5'h10: rom_data6_1 =  32'b10000000_00111111_11111100_00000000; 	//   *         ************         *
	5'h11: rom_data6_1 =  32'b10000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h12: rom_data6_1 =  32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h13: rom_data6_1 =  32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h14: rom_data6_1 =  32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h15: rom_data6_1 =  32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h16: rom_data6_1 =  32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h17: rom_data6_1 =  32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h18: rom_data6_1 =  32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h19: rom_data6_1 =  32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h1A: rom_data6_1 =  32'b10000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h1B: rom_data6_1 =  32'b10000000_00111111_11111100_00000000;	//   *         ************         *
	5'h1C: rom_data6_1 =  32'b10000000_00011111_11111000_00000000;	//   *          **********          *
	5'h1D: rom_data6_1 =  32'b10000000_00000000_00000000_00000000; 	//   *				    *
	5'h1E: rom_data6_1 =  32'b10000000_00000000_00000000_00000000; 	//   *				    *
	5'h1F: rom_data6_1 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr6_1 = pix_y[4:0] - NUM_y_t_1[4:0];
assign rom_col6_1 = pix_x[4:0] - NUM_x_l_1[4:0];

//------------------------------------//
// Number 7
wire [4:0] rom_addr7_1, rom_col7_1;
reg [31:0] rom_data7_1;

// number image ROM
always @*
case (rom_addr7_1)
	5'h0: rom_data7_1 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data7_1 =   32'b10000000_00000000_00000000_00000000;	//   *                              *
	5'h2: rom_data7_1 =   32'b10000000_00000000_00000000_00000000;	//   *                              *
	5'h3: rom_data7_1 =   32'b10000000_00011111_11111000_00000000;	//   *          **********          *
	5'h4: rom_data7_1 =   32'b10000000_00111111_11111100_00000000;	//   *         ************         *
	5'h5: rom_data7_1 =   32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h6: rom_data7_1 =   32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h7: rom_data7_1 =   32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h8: rom_data7_1 =   32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h9: rom_data7_1 =   32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'hA: rom_data7_1 =   32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'hB: rom_data7_1 =   32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'hC: rom_data7_1 =   32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'hD: rom_data7_1 =   32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'hE: rom_data7_1 =   32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'hF: rom_data7_1 =   32'b10000000_01000000_00000000_00000000;	//   *        *                     *
	5'h10: rom_data7_1 =  32'b10000000_01000000_00000000_00000000;	//   *        *                     *
	5'h11: rom_data7_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h12: rom_data7_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h13: rom_data7_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h14: rom_data7_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h15: rom_data7_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h16: rom_data7_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h17: rom_data7_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h18: rom_data7_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h19: rom_data7_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h1A: rom_data7_1 =  32'b10000000_01000000_00000000_00000000;	//   *        *                     *
	5'h1B: rom_data7_1 =  32'b10000000_00000000_00000000_00000000; 	//   *				    *
	5'h1C: rom_data7_1 =  32'b10000000_00000000_00000000_00000000; 	//   *				    *
	5'h1D: rom_data7_1 =  32'b10000000_00000000_00000000_00000000; 	//   *				    *
	5'h1E: rom_data7_1 =  32'b10000000_00000000_00000000_00000000; 	//   *				    *
	5'h1F: rom_data7_1 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr7_1 = pix_y[4:0] - NUM_y_t_1[4:0];
assign rom_col7_1 = pix_x[4:0] - NUM_x_l_1[4:0];

//------------------------------------//
// Number 8
wire [4:0] rom_addr8_1, rom_col8_1;
reg [31:0] rom_data8_1;

// number image ROM
always @*
case (rom_addr8_1)
	5'h0: rom_data8_1 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data8_1 =   32'b10000000_00000000_00000000_00000000;	//   *                              *
	5'h2: rom_data8_1 =   32'b10000000_00000000_00000000_00000000;	//   *                              *
	5'h3: rom_data8_1 =   32'b10000000_00011111_11111000_00000000;	//   *          **********          *
	5'h4: rom_data8_1 =   32'b10000000_00111111_11111100_00000000;	//   *         ************         *
	5'h5: rom_data8_1 =   32'b10000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h6: rom_data8_1 =   32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h7: rom_data8_1 =   32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h8: rom_data8_1 =   32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h9: rom_data8_1 =   32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hA: rom_data8_1 =   32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hB: rom_data8_1 =   32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hC: rom_data8_1 =   32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hD: rom_data8_1 =   32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hE: rom_data8_1 =   32'b10000000_01000000_00000010_00000000;	//   *        *            *        *
	5'hF: rom_data8_1 =   32'b10000000_00111111_11111100_00000000;	//   *         ************         *
	5'h10: rom_data8_1 =  32'b10000000_00111111_11111100_00000000; 	//   *         ************         *
	5'h11: rom_data8_1 =  32'b10000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h12: rom_data8_1 =  32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h13: rom_data8_1 =  32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h14: rom_data8_1 =  32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h15: rom_data8_1 =  32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h16: rom_data8_1 =  32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h17: rom_data8_1 =  32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h18: rom_data8_1 =  32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h19: rom_data8_1 =  32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h1A: rom_data8_1 =  32'b10000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h1B: rom_data8_1 =  32'b10000000_00111111_11111100_00000000;	//   *         ************         *
	5'h1C: rom_data8_1 =  32'b10000000_00011111_11111000_00000000;	//   *          **********          *
	5'h1D: rom_data8_1 =  32'b10000000_00000000_00000000_00000000; 	//   *				    *
	5'h1E: rom_data8_1 =  32'b10000000_00000000_00000000_00000000; 	//   *				    *
	5'h1F: rom_data8_1 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr8_1 = pix_y[4:0] - NUM_y_t_1[4:0];
assign rom_col8_1 = pix_x[4:0] - NUM_x_l_1[4:0];

//------------------------------------//
// Number 9
wire [4:0] rom_addr9_1, rom_col9_1;
reg [31:0] rom_data9_1;

// number image ROM
always @*
case (rom_addr9_1)
	5'h0: rom_data9_1 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data9_1 =   32'b10000000_00000000_00000000_00000000;	//   *                              *
	5'h2: rom_data9_1 =   32'b10000000_00000000_00000000_00000000;	//   *                              *
	5'h3: rom_data9_1 =   32'b10000000_00011111_11111000_00000000;	//   *          **********          *
	5'h4: rom_data9_1 =   32'b10000000_00111111_11111100_00000000;	//   *         ************         *
	5'h5: rom_data9_1 =   32'b10000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h6: rom_data9_1 =   32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h7: rom_data9_1 =   32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h8: rom_data9_1 =   32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h9: rom_data9_1 =   32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hA: rom_data9_1 =   32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hB: rom_data9_1 =   32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hC: rom_data9_1 =   32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hD: rom_data9_1 =   32'b10000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hE: rom_data9_1 =   32'b10000000_01000000_00000010_00000000;	//   *        *            *        *
	5'hF: rom_data9_1 =   32'b10000000_00111111_11111100_00000000;	//   *         ************         *
	5'h10: rom_data9_1 =  32'b10000000_00111111_11111100_00000000; 	//   *         ************         *
	5'h11: rom_data9_1 =  32'b10000000_01000000_00000000_00000000;	//   *        *                     *
	5'h12: rom_data9_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h13: rom_data9_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h14: rom_data9_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h15: rom_data9_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h16: rom_data9_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h17: rom_data9_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h18: rom_data9_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h19: rom_data9_1 =  32'b10000000_11000000_00000000_00000000;	//   *       **                     *
	5'h1A: rom_data9_1 =  32'b10000000_01000000_00000000_00000000;	//   *        *                     *
	5'h1B: rom_data9_1 =  32'b10000000_00000000_00000000_00000000; 	//   *				    *
	5'h1C: rom_data9_1 =  32'b10000000_00000000_00000000_00000000; 	//   *				    *
	5'h1D: rom_data9_1 =  32'b10000000_00000000_00000000_00000000; 	//   *				    *
	5'h1E: rom_data9_1 =  32'b10000000_00000000_00000000_00000000; 	//   *				    *
	5'h1F: rom_data9_1 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr9_1 = pix_y[4:0] - NUM_y_t_1[4:0];
assign rom_col9_1 = pix_x[4:0] - NUM_x_l_1[4:0];

always @(posedge clk) begin
	if (score[3:0] == 0)
	    rom_bit_1 = rom_data0_1[rom_col0_1];
	else if (score[3:0] == 1)
	    rom_bit_1 = rom_data1_1[rom_col1_1];
	else if (score[3:0] == 2)
	    rom_bit_1 = rom_data2_1[rom_col2_1];
	else if (score[3:0] == 3)
	    rom_bit_1 = rom_data3_1[rom_col3_1];
	else if (score[3:0] == 4)
	    rom_bit_1 = rom_data4_1[rom_col4_1];
	else if (score[3:0] == 5)
	    rom_bit_1 = rom_data5_1[rom_col5_1];
	else if (score[3:0] == 6)
	    rom_bit_1 = rom_data6_1[rom_col6_1];
	else if (score[3:0] == 7)
	    rom_bit_1 = rom_data7_1[rom_col7_1];
	else if (score[3:0] == 8)
	    rom_bit_1 = rom_data8_1[rom_col8_1];
	else if (score[3:0] == 9)
	    rom_bit_1 = rom_data9_1[rom_col9_1];
end


//-------------------------------------------------------------------------------------------------------------//
// Middle - Right Number

// number left, right boundary
wire [10:0] NUM_x_l_12 = 400;
wire [10:0] NUM_x_r_12 = NUM_x_l_12 + NUM_SIZE - 1;
// number top, bottom boundary 
wire [10:0] NUM_y_t_12 = 565; 
wire [10:0] NUM_y_b_12 = NUM_y_t_12 + NUM_SIZE - 1;
reg rom_bit_12;

//------------------------------------//
// Number 0
wire [4:0] rom_addr0_12, rom_col0_12;
reg [31:0] rom_data0_12;

// number image ROM
always @*
case (rom_addr0_12)
	5'h0: rom_data0_12 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data0_12 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h2: rom_data0_12 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h3: rom_data0_12 =   32'b00000000_00011111_11111000_00000000;	//   *          **********          *
	5'h4: rom_data0_12 =   32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h5: rom_data0_12 =   32'b00000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h6: rom_data0_12 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h7: rom_data0_12 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h8: rom_data0_12 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h9: rom_data0_12 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hA: rom_data0_12 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hB: rom_data0_12 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hC: rom_data0_12 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hD: rom_data0_12 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hE: rom_data0_12 =   32'b00000000_01000000_00000010_00000000;	//   *        *            *        *
	5'hF: rom_data0_12 =   32'b00000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h10: rom_data0_12 =  32'b00000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h11: rom_data0_12 =  32'b00000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h12: rom_data0_12 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h13: rom_data0_12 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h14: rom_data0_12 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h15: rom_data0_12 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h16: rom_data0_12 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h17: rom_data0_12 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h18: rom_data0_12 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h19: rom_data0_12 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h1A: rom_data0_12 =  32'b00000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h1B: rom_data0_12 =  32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h1C: rom_data0_12 =  32'b00000000_00011111_11111000_00000000;	//   *          **********          *
	5'h1D: rom_data0_12 =  32'b00000000_00000000_00000000_00000000; //   *				    *
	5'h1E: rom_data0_12 =  32'b00000000_00000000_00000000_00000000; //   *				    *
	5'h1F: rom_data0_12 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr0_12 = pix_y[4:0] - NUM_y_t_12[4:0];
assign rom_col0_12 = pix_x[4:0] - NUM_x_l_12[4:0];

//------------------------------------//
// Number 1
wire [4:0] rom_addr1_12, rom_col1_12;
reg [31:0] rom_data1_12;

// number image ROM
always @*
case (rom_addr1_12)
	5'h0: rom_data1_12 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data1_12 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h2: rom_data1_12 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h3: rom_data1_12 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h4: rom_data1_12 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h5: rom_data1_12 =   32'b00000000_01000000_00000000_00000000;	//   *        *                     *
	5'h6: rom_data1_12 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h7: rom_data1_12 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h8: rom_data1_12 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h9: rom_data1_12 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hA: rom_data1_12 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hB: rom_data1_12 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hC: rom_data1_12 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hD: rom_data1_12 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hE: rom_data1_12 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hF: rom_data1_12 =   32'b00000000_01000000_00000000_00000000;	//   *        *                     *
	5'h10: rom_data1_12 =  32'b00000000_01000000_00000000_00000000;	//   *        *                     *
	5'h11: rom_data1_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h12: rom_data1_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h13: rom_data1_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h14: rom_data1_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h15: rom_data1_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h16: rom_data1_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h17: rom_data1_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h18: rom_data1_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h19: rom_data1_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h1A: rom_data1_12 =  32'b00000000_01000000_00000000_00000000;	//   *        *                     *
	5'h1B: rom_data1_12 =  32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h1C: rom_data1_12 =  32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h1D: rom_data1_12 =  32'b00000000_00000000_00000000_00000000; //   *				    *
	5'h1E: rom_data1_12 =  32'b00000000_00000000_00000000_00000000; //   *				    *
	5'h1F: rom_data1_12 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr1_12 = pix_y[4:0] - NUM_y_t_12[4:0];
assign rom_col1_12 = pix_x[4:0] - NUM_x_l_12[4:0];

//------------------------------------//
// Number 2
wire [4:0] rom_addr2_12, rom_col2_12;
reg [31:0] rom_data2_12;

// number image ROM
always @*
case (rom_addr2_12)
	5'h0: rom_data2_12 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data2_12 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h2: rom_data2_12 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h3: rom_data2_12 =   32'b00000000_00011111_11111000_00000000;	//   *          **********          *
	5'h4: rom_data2_12 =   32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h5: rom_data2_12 =   32'b00000000_01000000_00000000_00000000;	//   *        *                     *
	5'h6: rom_data2_12 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h7: rom_data2_12 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h8: rom_data2_12 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h9: rom_data2_12 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hA: rom_data2_12 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hB: rom_data2_12 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hC: rom_data2_12 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hD: rom_data2_12 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hE: rom_data2_12 =   32'b00000000_01000000_00000000_00000000;	//   *        *                     *
	5'hF: rom_data2_12 =   32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h10: rom_data2_12 =  32'b00000000_00111111_11111100_00000000; //   *         ************         *
	5'h11: rom_data2_12 =  32'b00000000_00000000_00000010_00000000;	//   *                     *        *
	5'h12: rom_data2_12 =  32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'h13: rom_data2_12 =  32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'h14: rom_data2_12 =  32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'h15: rom_data2_12 =  32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'h16: rom_data2_12 =  32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'h17: rom_data2_12 =  32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'h18: rom_data2_12 =  32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'h19: rom_data2_12 =  32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'h1A: rom_data2_12 =  32'b00000000_00000000_00000010_00000000;	//   *                     *        *
	5'h1B: rom_data2_12 =  32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h1C: rom_data2_12 =  32'b00000000_00011111_11111000_00000000;	//   *          **********          *
	5'h1D: rom_data2_12 =  32'b00000000_00000000_00000000_00000000; //   *				    *
	5'h1E: rom_data2_12 =  32'b00000000_00000000_00000000_00000000; //   *				    *
	5'h1F: rom_data2_12 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr2_12 = pix_y[4:0] - NUM_y_t_12[4:0];
assign rom_col2_12 = pix_x[4:0] - NUM_x_l_12[4:0];

//------------------------------------//
// Number 3
wire [4:0] rom_addr3_12, rom_col3_12;
reg [31:0] rom_data3_12;

// number image ROM
always @*
case (rom_addr3_12)
	5'h0: rom_data3_12 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data3_12 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h2: rom_data3_12 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h3: rom_data3_12 =   32'b00000000_00011111_11111000_00000000;	//   *          **********          *
	5'h4: rom_data3_12 =   32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h5: rom_data3_12 =   32'b00000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h6: rom_data3_12 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h7: rom_data3_12 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h8: rom_data3_12 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h9: rom_data3_12 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hA: rom_data3_12 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hB: rom_data3_12 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hC: rom_data3_12 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hD: rom_data3_12 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hE: rom_data3_12 =   32'b00000000_01000000_00000000_00000000;	//   *        *                     *
	5'hF: rom_data3_12 =   32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h10: rom_data3_12 =  32'b00000000_00111111_11111100_00000000; //   *         ************         *
	5'h11: rom_data3_12 =  32'b00000000_01000000_00000000_00000000;	//   *        *                     *
	5'h12: rom_data3_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h13: rom_data3_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h14: rom_data3_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h15: rom_data3_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h16: rom_data3_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h17: rom_data3_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h18: rom_data3_12 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h19: rom_data3_12 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h1A: rom_data3_12 =  32'b00000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h1B: rom_data3_12 =  32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h1C: rom_data3_12 =  32'b00000000_00011111_11111000_00000000;	//   *          **********          *
	5'h1D: rom_data3_12 =  32'b00000000_00000000_00000000_00000000; //   *				    *
	5'h1E: rom_data3_12 =  32'b00000000_00000000_00000000_00000000; //   *				    *
	5'h1F: rom_data3_12 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr3_12 = pix_y[4:0] - NUM_y_t_12[4:0];
assign rom_col3_12 = pix_x[4:0] - NUM_x_l_12[4:0];

//------------------------------------//
// Number 4
wire [4:0] rom_addr4_12, rom_col4_12;
reg [31:0] rom_data4_12;

// number image ROM
always @*
case (rom_addr4_12)
	5'h0: rom_data4_12 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data4_12 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h2: rom_data4_12 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h3: rom_data4_12 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h4: rom_data4_12 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h5: rom_data4_12 =   32'b00000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h6: rom_data4_12 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h7: rom_data4_12 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h8: rom_data4_12 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h9: rom_data4_12 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hA: rom_data4_12 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hB: rom_data4_12 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hC: rom_data4_12 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hD: rom_data4_12 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hE: rom_data4_12 =   32'b00000000_01000000_00000010_00000000;	//   *        *            *        *
	5'hF: rom_data4_12 =   32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h10: rom_data4_12 =  32'b00000000_00111111_11111100_00000000; //   *         ************         *
	5'h11: rom_data4_12 =  32'b00000000_01000000_00000000_00000000;	//   *        *                     *
	5'h12: rom_data4_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h13: rom_data4_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h14: rom_data4_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h15: rom_data4_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h16: rom_data4_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h17: rom_data4_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h18: rom_data4_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h19: rom_data4_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h1A: rom_data4_12 =  32'b00000000_01000000_00000000_00000000;	//   *        *                     *
	5'h1B: rom_data4_12 =  32'b00000000_00000000_00000000_00000000; //   *				    *
	5'h1C: rom_data4_12 =  32'b00000000_00000000_00000000_00000000; //   *				    *
	5'h1D: rom_data4_12 =  32'b00000000_00000000_00000000_00000000; //   *				    *
	5'h1E: rom_data4_12 =  32'b00000000_00000000_00000000_00000000; //   *				    *
	5'h1F: rom_data4_12 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr4_12 = pix_y[4:0] - NUM_y_t_12[4:0];
assign rom_col4_12 = pix_x[4:0] - NUM_x_l_12[4:0];

//------------------------------------//
// Number 5
wire [4:0] rom_addr5_12, rom_col5_12;
reg [31:0] rom_data5_12;

// number image ROM
always @*
case (rom_addr5_12)
	5'h0: rom_data5_12 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data5_12 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h2: rom_data5_12 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h3: rom_data5_12 =   32'b00000000_00011111_11111000_00000000;	//   *          **********          *
	5'h4: rom_data5_12 =   32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h5: rom_data5_12 =   32'b00000000_00000000_00000010_00000000;	//   *                     *        *
	5'h6: rom_data5_12 =   32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'h7: rom_data5_12 =   32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'h8: rom_data5_12 =   32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'h9: rom_data5_12 =   32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'hA: rom_data5_12 =   32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'hB: rom_data5_12 =   32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'hC: rom_data5_12 =   32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'hD: rom_data5_12 =   32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'hE: rom_data5_12 =   32'b00000000_00000000_00000010_00000000;	//   *                     *        *
	5'hF: rom_data5_12 =   32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h10: rom_data5_12 =  32'b00000000_00111111_11111100_00000000; //   *         ************         *
	5'h11: rom_data5_12 =  32'b00000000_01000000_00000000_00000000;	//   *        *                     *
	5'h12: rom_data5_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h13: rom_data5_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h14: rom_data5_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h15: rom_data5_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h16: rom_data5_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h17: rom_data5_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h18: rom_data5_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h19: rom_data5_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h1A: rom_data5_12 =  32'b00000000_01000000_00000000_00000000;	//   *        *                     *
	5'h1B: rom_data5_12 =  32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h1C: rom_data5_12 =  32'b00000000_00011111_11111000_00000000;	//   *          **********          *
	5'h1D: rom_data5_12 =  32'b00000000_00000000_00000000_00000000; //   *				    *
	5'h1E: rom_data5_12 =  32'b00000000_00000000_00000000_00000000; //   *				    *
	5'h1F: rom_data5_12 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr5_12 = pix_y[4:0] - NUM_y_t_12[4:0];
assign rom_col5_12 = pix_x[4:0] - NUM_x_l_12[4:0];

//------------------------------------//
// Number 6
wire [4:0] rom_addr6_12, rom_col6_12;
reg [31:0] rom_data6_12;

// number image ROM
always @*
case (rom_addr6_12)
	5'h0: rom_data6_12 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data6_12 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h2: rom_data6_12 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h3: rom_data6_12 =   32'b00000000_00011111_11111000_00000000;	//   *          **********          *
	5'h4: rom_data6_12 =   32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h5: rom_data6_12 =   32'b00000000_00000000_00000010_00000000;	//   *                     *        *
	5'h6: rom_data6_12 =   32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'h7: rom_data6_12 =   32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'h8: rom_data6_12 =   32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'h9: rom_data6_12 =   32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'hA: rom_data6_12 =   32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'hB: rom_data6_12 =   32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'hC: rom_data6_12 =   32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'hD: rom_data6_12 =   32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'hE: rom_data6_12 =   32'b00000000_00000000_00000010_00000000;	//   *                     *        *
	5'hF: rom_data6_12 =   32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h10: rom_data6_12 =  32'b00000000_00111111_11111100_00000000; //   *         ************         *
	5'h11: rom_data6_12 =  32'b00000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h12: rom_data6_12 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h13: rom_data6_12 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h14: rom_data6_12 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h15: rom_data6_12 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h16: rom_data6_12 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h17: rom_data6_12 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h18: rom_data6_12 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h19: rom_data6_12 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h1A: rom_data6_12 =  32'b00000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h1B: rom_data6_12 =  32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h1C: rom_data6_12 =  32'b00000000_00011111_11111000_00000000;	//   *          **********          *
	5'h1D: rom_data6_12 =  32'b00000000_00000000_00000000_00000000; //   *				    *
	5'h1E: rom_data6_12 =  32'b00000000_00000000_00000000_00000000; //   *				    *
	5'h1F: rom_data6_12 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr6_12 = pix_y[4:0] - NUM_y_t_12[4:0];
assign rom_col6_12 = pix_x[4:0] - NUM_x_l_12[4:0];

//------------------------------------//
// Number 7
wire [4:0] rom_addr7_12, rom_col7_12;
reg [31:0] rom_data7_12;

// number image ROM
always @*
case (rom_addr7_12)
	5'h0: rom_data7_12 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data7_12 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h2: rom_data7_12 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h3: rom_data7_12 =   32'b00000000_00011111_11111000_00000000;	//   *          **********          *
	5'h4: rom_data7_12 =   32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h5: rom_data7_12 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h6: rom_data7_12 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h7: rom_data7_12 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h8: rom_data7_12 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h9: rom_data7_12 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hA: rom_data7_12 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hB: rom_data7_12 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hC: rom_data7_12 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hD: rom_data7_12 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hE: rom_data7_12 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hF: rom_data7_12 =   32'b00000000_01000000_00000000_00000000;	//   *        *                     *
	5'h10: rom_data7_12 =  32'b00000000_01000000_00000000_00000000;	//   *        *                     *
	5'h11: rom_data7_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h12: rom_data7_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h13: rom_data7_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h14: rom_data7_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h15: rom_data7_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h16: rom_data7_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h17: rom_data7_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h18: rom_data7_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h19: rom_data7_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h1A: rom_data7_12 =  32'b00000000_01000000_00000000_00000000;	//   *        *                     *
	5'h1B: rom_data7_12 =  32'b00000000_00000000_00000000_00000000; //   *				    *
	5'h1C: rom_data7_12 =  32'b00000000_00000000_00000000_00000000; //   *				    *
	5'h1D: rom_data7_12 =  32'b00000000_00000000_00000000_00000000; //   *				    *
	5'h1E: rom_data7_12 =  32'b00000000_00000000_00000000_00000000; //   *				    *
	5'h1F: rom_data7_12 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr7_12 = pix_y[4:0] - NUM_y_t_12[4:0];
assign rom_col7_12 = pix_x[4:0] - NUM_x_l_12[4:0];

//------------------------------------//
// Number 8
wire [4:0] rom_addr8_12, rom_col8_12;
reg [31:0] rom_data8_12;

// number image ROM
always @*
case (rom_addr8_12)
	5'h0: rom_data8_12 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data8_12 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h2: rom_data8_12 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h3: rom_data8_12 =   32'b00000000_00011111_11111000_00000000;	//   *          **********          *
	5'h4: rom_data8_12 =   32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h5: rom_data8_12 =   32'b00000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h6: rom_data8_12 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h7: rom_data8_12 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h8: rom_data8_12 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h9: rom_data8_12 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hA: rom_data8_12 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hB: rom_data8_12 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hC: rom_data8_12 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hD: rom_data8_12 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hE: rom_data8_12 =   32'b00000000_01000000_00000010_00000000;	//   *        *            *        *
	5'hF: rom_data8_12 =   32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h10: rom_data8_12 =  32'b00000000_00111111_11111100_00000000; //   *         ************         *
	5'h11: rom_data8_12 =  32'b00000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h12: rom_data8_12 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h13: rom_data8_12 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h14: rom_data8_12 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h15: rom_data8_12 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h16: rom_data8_12 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h17: rom_data8_12 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h18: rom_data8_12 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h19: rom_data8_12 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h1A: rom_data8_12 =  32'b00000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h1B: rom_data8_12 =  32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h1C: rom_data8_12 =  32'b00000000_00011111_11111000_00000000;	//   *          **********          *
	5'h1D: rom_data8_12 =  32'b00000000_00000000_00000000_00000000; //   *				    *
	5'h1E: rom_data8_12 =  32'b00000000_00000000_00000000_00000000; //   *				    *
	5'h1F: rom_data8_12 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr8_12 = pix_y[4:0] - NUM_y_t_12[4:0];
assign rom_col8_12 = pix_x[4:0] - NUM_x_l_12[4:0];

//------------------------------------//
// Number 9
wire [4:0] rom_addr9_12, rom_col9_12;
reg [31:0] rom_data9_12;

// number image ROM
always @*
case (rom_addr9_12)
	5'h0: rom_data9_12 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data9_12 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h2: rom_data9_12 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h3: rom_data9_12 =   32'b00000000_00011111_11111000_00000000;	//   *          **********          *
	5'h4: rom_data9_12 =   32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h5: rom_data9_12 =   32'b00000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h6: rom_data9_12 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h7: rom_data9_12 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h8: rom_data9_12 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h9: rom_data9_12 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hA: rom_data9_12 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hB: rom_data9_12 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hC: rom_data9_12 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hD: rom_data9_12 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hE: rom_data9_12 =   32'b00000000_01000000_00000010_00000000;	//   *        *            *        *
	5'hF: rom_data9_12 =   32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h10: rom_data9_12 =  32'b00000000_00111111_11111100_00000000; //   *         ************         *
	5'h11: rom_data9_12 =  32'b00000000_01000000_00000000_00000000;	//   *        *                     *
	5'h12: rom_data9_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h13: rom_data9_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h14: rom_data9_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h15: rom_data9_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h16: rom_data9_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h17: rom_data9_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h18: rom_data9_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h19: rom_data9_12 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h1A: rom_data9_12 =  32'b00000000_01000000_00000000_00000000;	//   *        *                     *
	5'h1B: rom_data9_12 =  32'b00000000_00000000_00000000_00000000; //   *				    *
	5'h1C: rom_data9_12 =  32'b00000000_00000000_00000000_00000000; //   *				    *
	5'h1D: rom_data9_12 =  32'b00000000_00000000_00000000_00000000; //   *				    *
	5'h1E: rom_data9_12 =  32'b00000000_00000000_00000000_00000000; //   *				    *
	5'h1F: rom_data9_12 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr9_12 = pix_y[4:0] - NUM_y_t_12[4:0];
assign rom_col9_12 = pix_x[4:0] - NUM_x_l_12[4:0];

always @(posedge clk) begin
	if (score[7:4] == 0)
	    rom_bit_12 = rom_data0_12[rom_col0_12];
	else if (score[7:4] == 1)
	    rom_bit_12 = rom_data1_12[rom_col1_12];
	else if (score[7:4] == 2)
	    rom_bit_12 = rom_data2_12[rom_col2_12];
	else if (score[7:4] == 3)
	    rom_bit_12 = rom_data3_12[rom_col3_12];
	else if (score[7:4] == 4)
	    rom_bit_12 = rom_data4_12[rom_col4_12];
	else if (score[7:4] == 5)
	    rom_bit_12 = rom_data5_12[rom_col5_12];
	else if (score[7:4] == 6)
	    rom_bit_12 = rom_data6_12[rom_col6_12];
	else if (score[7:4] == 7)
	    rom_bit_12 = rom_data7_12[rom_col7_12];
	else if (score[7:4] == 8)
	    rom_bit_12 = rom_data8_12[rom_col8_12];
	else if (score[7:4] == 9)
	    rom_bit_12 = rom_data9_12[rom_col9_12];
end


//-------------------------------------------------------------------------------------------------------------//
// Middle - Left Number

// number left, right boundary
wire [10:0] NUM_x_l_123 = 368;
wire [10:0] NUM_x_r_123 = NUM_x_l_123 + NUM_SIZE - 1;
// number top, bottom boundary 
wire [10:0] NUM_y_t_123 = 565; 
wire [10:0] NUM_y_b_123 = NUM_y_t_123 + NUM_SIZE - 1;
reg rom_bit_123;

//------------------------------------//
// Number 0
wire [4:0] rom_addr0_123, rom_col0_123;
reg [31:0] rom_data0_123;

// number image ROM
always @*
case (rom_addr0_123)
	5'h0: rom_data0_123 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data0_123 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h2: rom_data0_123 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h3: rom_data0_123 =   32'b00000000_00011111_11111000_00000000;	//   *          **********          *
	5'h4: rom_data0_123 =   32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h5: rom_data0_123 =   32'b00000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h6: rom_data0_123 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h7: rom_data0_123 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h8: rom_data0_123 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h9: rom_data0_123 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hA: rom_data0_123 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hB: rom_data0_123 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hC: rom_data0_123 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hD: rom_data0_123 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hE: rom_data0_123 =   32'b00000000_01000000_00000010_00000000;	//   *        *            *        *
	5'hF: rom_data0_123 =   32'b00000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h10: rom_data0_123 =  32'b00000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h11: rom_data0_123 =  32'b00000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h12: rom_data0_123 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h13: rom_data0_123 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h14: rom_data0_123 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h15: rom_data0_123 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h16: rom_data0_123 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h17: rom_data0_123 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h18: rom_data0_123 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h19: rom_data0_123 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h1A: rom_data0_123 =  32'b00000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h1B: rom_data0_123 =  32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h1C: rom_data0_123 =  32'b00000000_00011111_11111000_00000000;	//   *          **********          *
	5'h1D: rom_data0_123 =  32'b00000000_00000000_00000000_00000000; 	//   *				    *
	5'h1E: rom_data0_123 =  32'b00000000_00000000_00000000_00000000; 	//   *				    *
	5'h1F: rom_data0_123 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr0_123 = pix_y[4:0] - NUM_y_t_123[4:0];
assign rom_col0_123 = pix_x[4:0] - NUM_x_l_123[4:0];

//------------------------------------//
// Number 1
wire [4:0] rom_addr1_123, rom_col1_123;
reg [31:0] rom_data1_123;

// number image ROM
always @*
case (rom_addr1_123)
	5'h0: rom_data1_123 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data1_123 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h2: rom_data1_123 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h3: rom_data1_123 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h4: rom_data1_123 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h5: rom_data1_123 =   32'b00000000_01000000_00000000_00000000;	//   *        *                     *
	5'h6: rom_data1_123 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h7: rom_data1_123 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h8: rom_data1_123 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h9: rom_data1_123 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hA: rom_data1_123 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hB: rom_data1_123 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hC: rom_data1_123 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hD: rom_data1_123 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hE: rom_data1_123 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hF: rom_data1_123 =   32'b00000000_01000000_00000000_00000000;	//   *        *                     *
	5'h10: rom_data1_123 =  32'b00000000_01000000_00000000_00000000;	//   *        *                     *
	5'h11: rom_data1_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h12: rom_data1_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h13: rom_data1_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h14: rom_data1_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h15: rom_data1_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h16: rom_data1_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h17: rom_data1_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h18: rom_data1_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h19: rom_data1_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h1A: rom_data1_123 =  32'b00000000_01000000_00000000_00000000;	//   *        *                     *
	5'h1B: rom_data1_123 =  32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h1C: rom_data1_123 =  32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h1D: rom_data1_123 =  32'b00000000_00000000_00000000_00000000; 	//   *				    *
	5'h1E: rom_data1_123 =  32'b00000000_00000000_00000000_00000000; 	//   *				    *
	5'h1F: rom_data1_123 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr1_123 = pix_y[4:0] - NUM_y_t_123[4:0];
assign rom_col1_123 = pix_x[4:0] - NUM_x_l_123[4:0];

//------------------------------------//
// Number 2
wire [4:0] rom_addr2_123, rom_col2_123;
reg [31:0] rom_data2_123;

// number image ROM
always @*
case (rom_addr2_123)
	5'h0: rom_data2_123 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data2_123 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h2: rom_data2_123 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h3: rom_data2_123 =   32'b00000000_00011111_11111000_00000000;	//   *          **********          *
	5'h4: rom_data2_123 =   32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h5: rom_data2_123 =   32'b00000000_01000000_00000000_00000000;	//   *        *                     *
	5'h6: rom_data2_123 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h7: rom_data2_123 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h8: rom_data2_123 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h9: rom_data2_123 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hA: rom_data2_123 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hB: rom_data2_123 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hC: rom_data2_123 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hD: rom_data2_123 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hE: rom_data2_123 =   32'b00000000_01000000_00000000_00000000;	//   *        *                     *
	5'hF: rom_data2_123 =   32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h10: rom_data2_123 =  32'b00000000_00111111_11111100_00000000; 	//   *         ************         *
	5'h11: rom_data2_123 =  32'b00000000_00000000_00000010_00000000;	//   *                     *        *
	5'h12: rom_data2_123 =  32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'h13: rom_data2_123 =  32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'h14: rom_data2_123 =  32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'h15: rom_data2_123 =  32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'h16: rom_data2_123 =  32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'h17: rom_data2_123 =  32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'h18: rom_data2_123 =  32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'h19: rom_data2_123 =  32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'h1A: rom_data2_123 =  32'b00000000_00000000_00000010_00000000;	//   *                     *        *
	5'h1B: rom_data2_123 =  32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h1C: rom_data2_123 =  32'b00000000_00011111_11111000_00000000;	//   *          **********          *
	5'h1D: rom_data2_123 =  32'b00000000_00000000_00000000_00000000; 	//   *				    *
	5'h1E: rom_data2_123 =  32'b00000000_00000000_00000000_00000000; 	//   *				    *
	5'h1F: rom_data2_123 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr2_123 = pix_y[4:0] - NUM_y_t_123[4:0];
assign rom_col2_123 = pix_x[4:0] - NUM_x_l_123[4:0];

//------------------------------------//
// Number 3
wire [4:0] rom_addr3_123, rom_col3_123;
reg [31:0] rom_data3_123;

// number image ROM
always @*
case (rom_addr3_123)
	5'h0: rom_data3_123 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data3_123 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h2: rom_data3_123 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h3: rom_data3_123 =   32'b00000000_00011111_11111000_00000000;	//   *          **********          *
	5'h4: rom_data3_123 =   32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h5: rom_data3_123 =   32'b00000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h6: rom_data3_123 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h7: rom_data3_123 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h8: rom_data3_123 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h9: rom_data3_123 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hA: rom_data3_123 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hB: rom_data3_123 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hC: rom_data3_123 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hD: rom_data3_123 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hE: rom_data3_123 =   32'b00000000_01000000_00000000_00000000;	//   *        *                     *
	5'hF: rom_data3_123 =   32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h10: rom_data3_123 =  32'b00000000_00111111_11111100_00000000; 	//   *         ************         *
	5'h11: rom_data3_123 =  32'b00000000_01000000_00000000_00000000;	//   *        *                     *
	5'h12: rom_data3_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h13: rom_data3_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h14: rom_data3_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h15: rom_data3_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h16: rom_data3_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h17: rom_data3_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h18: rom_data3_123 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h19: rom_data3_123 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h1A: rom_data3_123 =  32'b00000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h1B: rom_data3_123 =  32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h1C: rom_data3_123 =  32'b00000000_00011111_11111000_00000000;	//   *          **********          *
	5'h1D: rom_data3_123 =  32'b00000000_00000000_00000000_00000000; 	//   *				    *
	5'h1E: rom_data3_123 =  32'b00000000_00000000_00000000_00000000; 	//   *				    *
	5'h1F: rom_data3_123 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr3_123 = pix_y[4:0] - NUM_y_t_123[4:0];
assign rom_col3_123 = pix_x[4:0] - NUM_x_l_123[4:0];

//------------------------------------//
// Number 4
wire [4:0] rom_addr4_123, rom_col4_123;
reg [31:0] rom_data4_123;

// number image ROM
always @*
case (rom_addr4_123)
	5'h0: rom_data4_123 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data4_123 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h2: rom_data4_123 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h3: rom_data4_123 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h4: rom_data4_123 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h5: rom_data4_123 =   32'b00000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h6: rom_data4_123 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h7: rom_data4_123 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h8: rom_data4_123 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h9: rom_data4_123 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hA: rom_data4_123 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hB: rom_data4_123 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hC: rom_data4_123 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hD: rom_data4_123 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hE: rom_data4_123 =   32'b00000000_01000000_00000010_00000000;	//   *        *            *        *
	5'hF: rom_data4_123 =   32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h10: rom_data4_123 =  32'b00000000_00111111_11111100_00000000; 	//   *         ************         *
	5'h11: rom_data4_123 =  32'b00000000_01000000_00000000_00000000;	//   *        *                     *
	5'h12: rom_data4_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h13: rom_data4_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h14: rom_data4_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h15: rom_data4_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h16: rom_data4_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h17: rom_data4_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h18: rom_data4_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h19: rom_data4_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h1A: rom_data4_123 =  32'b00000000_01000000_00000000_00000000;	//   *        *                     *
	5'h1B: rom_data4_123 =  32'b00000000_00000000_00000000_00000000; 	//   *				    *
	5'h1C: rom_data4_123 =  32'b00000000_00000000_00000000_00000000; 	//   *				    *
	5'h1D: rom_data4_123 =  32'b00000000_00000000_00000000_00000000; 	//   *				    *
	5'h1E: rom_data4_123 =  32'b00000000_00000000_00000000_00000000; 	//   *				    *
	5'h1F: rom_data4_123 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr4_123 = pix_y[4:0] - NUM_y_t_123[4:0];
assign rom_col4_123 = pix_x[4:0] - NUM_x_l_123[4:0];

//------------------------------------//
// Number 5
wire [4:0] rom_addr5_123, rom_col5_123;
reg [31:0] rom_data5_123;

// number image ROM
always @*
case (rom_addr5_123)
	5'h0: rom_data5_123 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data5_123 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h2: rom_data5_123 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h3: rom_data5_123 =   32'b00000000_00011111_11111000_00000000;	//   *          **********          *
	5'h4: rom_data5_123 =   32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h5: rom_data5_123 =   32'b00000000_00000000_00000010_00000000;	//   *                     *        *
	5'h6: rom_data5_123 =   32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'h7: rom_data5_123 =   32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'h8: rom_data5_123 =   32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'h9: rom_data5_123 =   32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'hA: rom_data5_123 =   32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'hB: rom_data5_123 =   32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'hC: rom_data5_123 =   32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'hD: rom_data5_123 =   32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'hE: rom_data5_123 =   32'b00000000_00000000_00000010_00000000;	//   *                     *        *
	5'hF: rom_data5_123 =   32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h10: rom_data5_123 =  32'b00000000_00111111_11111100_00000000; 	//   *         ************         *
	5'h11: rom_data5_123 =  32'b00000000_01000000_00000000_00000000;	//   *        *                     *
	5'h12: rom_data5_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h13: rom_data5_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h14: rom_data5_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h15: rom_data5_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h16: rom_data5_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h17: rom_data5_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h18: rom_data5_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h19: rom_data5_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h1A: rom_data5_123 =  32'b00000000_01000000_00000000_00000000;	//   *        *                     *
	5'h1B: rom_data5_123 =  32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h1C: rom_data5_123 =  32'b00000000_00011111_11111000_00000000;	//   *          **********          *
	5'h1D: rom_data5_123 =  32'b00000000_00000000_00000000_00000000; 	//   *				    *
	5'h1E: rom_data5_123 =  32'b00000000_00000000_00000000_00000000; 	//   *				    *
	5'h1F: rom_data5_123 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr5_123 = pix_y[4:0] - NUM_y_t_123[4:0];
assign rom_col5_123 = pix_x[4:0] - NUM_x_l_123[4:0];

//------------------------------------//
// Number 6
wire [4:0] rom_addr6_123, rom_col6_123;
reg [31:0] rom_data6_123;

// number image ROM
always @*
case (rom_addr6_123)
	5'h0: rom_data6_123 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data6_123 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h2: rom_data6_123 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h3: rom_data6_123 =   32'b00000000_00011111_11111000_00000000;	//   *          **********          *
	5'h4: rom_data6_123 =   32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h5: rom_data6_123 =   32'b00000000_00000000_00000010_00000000;	//   *                     *        *
	5'h6: rom_data6_123 =   32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'h7: rom_data6_123 =   32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'h8: rom_data6_123 =   32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'h9: rom_data6_123 =   32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'hA: rom_data6_123 =   32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'hB: rom_data6_123 =   32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'hC: rom_data6_123 =   32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'hD: rom_data6_123 =   32'b00000000_00000000_00000011_00000000;	//   *                     **       *
	5'hE: rom_data6_123 =   32'b00000000_00000000_00000010_00000000;	//   *                     *        *
	5'hF: rom_data6_123 =   32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h10: rom_data6_123 =  32'b00000000_00111111_11111100_00000000; 	//   *         ************         *
	5'h11: rom_data6_123 =  32'b00000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h12: rom_data6_123 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h13: rom_data6_123 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h14: rom_data6_123 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h15: rom_data6_123 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h16: rom_data6_123 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h17: rom_data6_123 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h18: rom_data6_123 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h19: rom_data6_123 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h1A: rom_data6_123 =  32'b00000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h1B: rom_data6_123 =  32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h1C: rom_data6_123 =  32'b00000000_00011111_11111000_00000000;	//   *          **********          *
	5'h1D: rom_data6_123 =  32'b00000000_00000000_00000000_00000000; 	//   *				    *
	5'h1E: rom_data6_123 =  32'b00000000_00000000_00000000_00000000; 	//   *				    *
	5'h1F: rom_data6_123 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr6_123 = pix_y[4:0] - NUM_y_t_123[4:0];
assign rom_col6_123 = pix_x[4:0] - NUM_x_l_123[4:0];

//------------------------------------//
// Number 7
wire [4:0] rom_addr7_123, rom_col7_123;
reg [31:0] rom_data7_123;

// number image ROM
always @*
case (rom_addr7_123)
	5'h0: rom_data7_123 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data7_123 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h2: rom_data7_123 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h3: rom_data7_123 =   32'b00000000_00011111_11111000_00000000;	//   *          **********          *
	5'h4: rom_data7_123 =   32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h5: rom_data7_123 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h6: rom_data7_123 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h7: rom_data7_123 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h8: rom_data7_123 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h9: rom_data7_123 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hA: rom_data7_123 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hB: rom_data7_123 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hC: rom_data7_123 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hD: rom_data7_123 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hE: rom_data7_123 =   32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'hF: rom_data7_123 =   32'b00000000_01000000_00000000_00000000;	//   *        *                     *
	5'h10: rom_data7_123 =  32'b00000000_01000000_00000000_00000000;	//   *        *                     *
	5'h11: rom_data7_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h12: rom_data7_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h13: rom_data7_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h14: rom_data7_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h15: rom_data7_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h16: rom_data7_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h17: rom_data7_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h18: rom_data7_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h19: rom_data7_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h1A: rom_data7_123 =  32'b00000000_01000000_00000000_00000000;	//   *        *                     *
	5'h1B: rom_data7_123 =  32'b00000000_00000000_00000000_00000000; 	//   *				    *
	5'h1C: rom_data7_123 =  32'b00000000_00000000_00000000_00000000; 	//   *				    *
	5'h1D: rom_data7_123 =  32'b00000000_00000000_00000000_00000000; 	//   *				    *
	5'h1E: rom_data7_123 =  32'b00000000_00000000_00000000_00000000; 	//   *				    *
	5'h1F: rom_data7_123 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr7_123 = pix_y[4:0] - NUM_y_t_123[4:0];
assign rom_col7_123 = pix_x[4:0] - NUM_x_l_123[4:0];

//------------------------------------//
// Number 8
wire [4:0] rom_addr8_123, rom_col8_123;
reg [31:0] rom_data8_123;

// number image ROM
always @*
case (rom_addr8_123)
	5'h0: rom_data8_123 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data8_123 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h2: rom_data8_123 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h3: rom_data8_123 =   32'b00000000_00011111_11111000_00000000;	//   *          **********          *
	5'h4: rom_data8_123 =   32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h5: rom_data8_123 =   32'b00000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h6: rom_data8_123 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h7: rom_data8_123 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h8: rom_data8_123 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h9: rom_data8_123 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hA: rom_data8_123 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hB: rom_data8_123 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hC: rom_data8_123 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hD: rom_data8_123 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hE: rom_data8_123 =   32'b00000000_01000000_00000010_00000000;	//   *        *            *        *
	5'hF: rom_data8_123 =   32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h10: rom_data8_123 =  32'b00000000_00111111_11111100_00000000; 	//   *         ************         *
	5'h11: rom_data8_123 =  32'b00000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h12: rom_data8_123 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h13: rom_data8_123 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h14: rom_data8_123 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h15: rom_data8_123 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h16: rom_data8_123 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h17: rom_data8_123 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h18: rom_data8_123 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h19: rom_data8_123 =  32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h1A: rom_data8_123 =  32'b00000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h1B: rom_data8_123 =  32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h1C: rom_data8_123 =  32'b00000000_00011111_11111000_00000000;	//   *          **********          *
	5'h1D: rom_data8_123 =  32'b00000000_00000000_00000000_00000000; 	//   *				    *
	5'h1E: rom_data8_123 =  32'b00000000_00000000_00000000_00000000; 	//   *				    *
	5'h1F: rom_data8_123 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr8_123 = pix_y[4:0] - NUM_y_t_123[4:0];
assign rom_col8_123 = pix_x[4:0] - NUM_x_l_123[4:0];

//------------------------------------//
// Number 9
wire [4:0] rom_addr9_123, rom_col9_123;
reg [31:0] rom_data9_123;

// number image ROM
always @*
case (rom_addr9_123)
	5'h0: rom_data9_123 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data9_123 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h2: rom_data9_123 =   32'b00000000_00000000_00000000_00000000;	//   *                              *
	5'h3: rom_data9_123 =   32'b00000000_00011111_11111000_00000000;	//   *          **********          *
	5'h4: rom_data9_123 =   32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h5: rom_data9_123 =   32'b00000000_01000000_00000010_00000000;	//   *        *            *        *
	5'h6: rom_data9_123 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h7: rom_data9_123 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h8: rom_data9_123 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'h9: rom_data9_123 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hA: rom_data9_123 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hB: rom_data9_123 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hC: rom_data9_123 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hD: rom_data9_123 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hE: rom_data9_123 =   32'b00000000_01000000_00000010_00000000;	//   *        *            *        *
	5'hF: rom_data9_123 =   32'b00000000_00111111_11111100_00000000;	//   *         ************         *
	5'h10: rom_data9_123 =  32'b00000000_00111111_11111100_00000000; 	//   *         ************         *
	5'h11: rom_data9_123 =  32'b00000000_01000000_00000000_00000000;	//   *        *                     *
	5'h12: rom_data9_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h13: rom_data9_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h14: rom_data9_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h15: rom_data9_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h16: rom_data9_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h17: rom_data9_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h18: rom_data9_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h19: rom_data9_123 =  32'b00000000_11000000_00000000_00000000;	//   *       **                     *
	5'h1A: rom_data9_123 =  32'b00000000_01000000_00000000_00000000;	//   *        *                     *
	5'h1B: rom_data9_123 =  32'b00000000_00000000_00000000_00000000; 	//   *				    *
	5'h1C: rom_data9_123 =  32'b00000000_00000000_00000000_00000000; 	//   *				    *
	5'h1D: rom_data9_123 =  32'b00000000_00000000_00000000_00000000; 	//   *				    *
	5'h1E: rom_data9_123 =  32'b00000000_00000000_00000000_00000000; 	//   *				    *
	5'h1F: rom_data9_123 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr9_123 = pix_y[4:0] - NUM_y_t_123[4:0];
assign rom_col9_123 = pix_x[4:0] - NUM_x_l_123[4:0];

always @(posedge clk) begin
	if (score[11:8] == 0)
	    rom_bit_123 = rom_data0_123[rom_col0_123];
	else if (score[11:8] == 1)
	    rom_bit_123 = rom_data1_123[rom_col1_123];
	else if (score[11:8] == 2)
	    rom_bit_123 = rom_data2_123[rom_col2_123];
	else if (score[11:8] == 3)
	    rom_bit_123 = rom_data3_123[rom_col3_123];
	else if (score[11:8] == 4)
	    rom_bit_123 = rom_data4_123[rom_col4_123];
	else if (score[11:8] == 5)
	    rom_bit_123 = rom_data5_123[rom_col5_123];
	else if (score[11:8] == 6)
	    rom_bit_123 = rom_data6_123[rom_col6_123];
	else if (score[11:8] == 7)
	    rom_bit_123 = rom_data7_123[rom_col7_123];
	else if (score[11:8] == 8)
	    rom_bit_123 = rom_data8_123[rom_col8_123];
	else if (score[11:8] == 9)
	    rom_bit_123 = rom_data9_123[rom_col9_123];
end

//-------------------------------------------------------------------------------------------------------------//
// Left Number

// number left, right boundary
wire [10:0] NUM_x_l_1234 = 336;
wire [10:0] NUM_x_r_1234 = NUM_x_l_1234 + NUM_SIZE - 1;
// number top, bottom boundary 
wire [10:0] NUM_y_t_1234 = 565; 
wire [10:0] NUM_y_b_1234 = NUM_y_t_1234 + NUM_SIZE - 1;
reg rom_bit_1234;

//------------------------------------//
// Number 0
wire [4:0] rom_addr0_1234, rom_col0_1234;
reg [31:0] rom_data0_1234;

// number image ROM
always @*
case (rom_addr0_1234)
	5'h0: rom_data0_1234 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data0_1234 =   32'b00000000_00000000_00000000_00000001;	//   *                              *
	5'h2: rom_data0_1234 =   32'b00000000_00000000_00000000_00000001;	//   *                              *
	5'h3: rom_data0_1234 =   32'b00000000_00011111_11111000_00000001;	//   *          **********          *
	5'h4: rom_data0_1234 =   32'b00000000_00111111_11111100_00000001;	//   *         ************         *
	5'h5: rom_data0_1234 =   32'b00000000_01000000_00000010_00000001;	//   *        *            *        *
	5'h6: rom_data0_1234 =   32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h7: rom_data0_1234 =   32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h8: rom_data0_1234 =   32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h9: rom_data0_1234 =   32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'hA: rom_data0_1234 =   32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'hB: rom_data0_1234 =   32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'hC: rom_data0_1234 =   32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'hD: rom_data0_1234 =   32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'hE: rom_data0_1234 =   32'b00000000_01000000_00000010_00000001;	//   *        *            *        *
	5'hF: rom_data0_1234 =   32'b00000000_01000000_00000010_00000001;	//   *        *            *        *
	5'h10: rom_data0_1234 =  32'b00000000_01000000_00000010_00000001;	//   *        *            *        *
	5'h11: rom_data0_1234 =  32'b00000000_01000000_00000010_00000001;	//   *        *            *        *
	5'h12: rom_data0_1234 =  32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h13: rom_data0_1234 =  32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h14: rom_data0_1234 =  32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h15: rom_data0_1234 =  32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h16: rom_data0_1234 =  32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h17: rom_data0_1234 =  32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h18: rom_data0_1234 =  32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h19: rom_data0_1234 =  32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h1A: rom_data0_1234 =  32'b00000000_01000000_00000010_00000001;	//   *        *            *        *
	5'h1B: rom_data0_1234 =  32'b00000000_00111111_11111100_00000001;	//   *         ************         *
	5'h1C: rom_data0_1234 =  32'b00000000_00011111_11111000_00000001;	//   *          **********          *
	5'h1D: rom_data0_1234 =  32'b00000000_00000000_00000000_00000001; 	//   *				    *
	5'h1E: rom_data0_1234 =  32'b00000000_00000000_00000000_00000001; 	//   *				    *
	5'h1F: rom_data0_1234 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr0_1234 = pix_y[4:0] - NUM_y_t_1234[4:0];
assign rom_col0_1234 = pix_x[4:0] - NUM_x_l_1234[4:0];

//------------------------------------//
// Number 1
wire [4:0] rom_addr1_1234, rom_col1_1234;
reg [31:0] rom_data1_1234;

// number image ROM
always @*
case (rom_addr1_1234)
	5'h0: rom_data1_1234 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data1_1234 =   32'b00000000_00000000_00000000_00000001;	//   *                              *
	5'h2: rom_data1_1234 =   32'b00000000_00000000_00000000_00000001;	//   *                              *
	5'h3: rom_data1_1234 =   32'b00000000_00000000_00000000_00000001;	//   *                              *
	5'h4: rom_data1_1234 =   32'b00000000_00000000_00000000_00000001;	//   *                              *
	5'h5: rom_data1_1234 =   32'b00000000_01000000_00000000_00000001;	//   *        *                     *
	5'h6: rom_data1_1234 =   32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h7: rom_data1_1234 =   32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h8: rom_data1_1234 =   32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h9: rom_data1_1234 =   32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'hA: rom_data1_1234 =   32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'hB: rom_data1_1234 =   32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'hC: rom_data1_1234 =   32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'hD: rom_data1_1234 =   32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'hE: rom_data1_1234 =   32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'hF: rom_data1_1234 =   32'b00000000_01000000_00000000_00000001;	//   *        *                     *
	5'h10: rom_data1_1234 =  32'b00000000_01000000_00000000_00000001;	//   *        *                     *
	5'h11: rom_data1_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h12: rom_data1_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h13: rom_data1_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h14: rom_data1_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h15: rom_data1_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h16: rom_data1_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h17: rom_data1_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h18: rom_data1_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h19: rom_data1_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h1A: rom_data1_1234 =  32'b00000000_01000000_00000000_00000001;	//   *        *                     *
	5'h1B: rom_data1_1234 =  32'b00000000_00000000_00000000_00000001;	//   *                              *
	5'h1C: rom_data1_1234 =  32'b00000000_00000000_00000000_00000001;	//   *                              *
	5'h1D: rom_data1_1234 =  32'b00000000_00000000_00000000_00000001; 	//   *				    *
	5'h1E: rom_data1_1234 =  32'b00000000_00000000_00000000_00000001; 	//   *				    *
	5'h1F: rom_data1_1234 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr1_1234 = pix_y[4:0] - NUM_y_t_1234[4:0];
assign rom_col1_1234 = pix_x[4:0] - NUM_x_l_1234[4:0];

//------------------------------------//
// Number 2
wire [4:0] rom_addr2_1234, rom_col2_1234;
reg [31:0] rom_data2_1234;

// number image ROM
always @*
case (rom_addr2_1234)
	5'h0: rom_data2_1234 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data2_1234 =   32'b00000000_00000000_00000000_00000001;	//   *                              *
	5'h2: rom_data2_1234 =   32'b00000000_00000000_00000000_00000001;	//   *                              *
	5'h3: rom_data2_1234 =   32'b00000000_00011111_11111000_00000001;	//   *          **********          *
	5'h4: rom_data2_1234 =   32'b00000000_00111111_11111100_00000001;	//   *         ************         *
	5'h5: rom_data2_1234 =   32'b00000000_01000000_00000000_00000001;	//   *        *                     *
	5'h6: rom_data2_1234 =   32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h7: rom_data2_1234 =   32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h8: rom_data2_1234 =   32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h9: rom_data2_1234 =   32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'hA: rom_data2_1234 =   32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'hB: rom_data2_1234 =   32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'hC: rom_data2_1234 =   32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'hD: rom_data2_1234 =   32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'hE: rom_data2_1234 =   32'b00000000_01000000_00000000_00000001;	//   *        *                     *
	5'hF: rom_data2_1234 =   32'b00000000_00111111_11111100_00000001;	//   *         ************         *
	5'h10: rom_data2_1234 =  32'b00000000_00111111_11111100_00000001; 	//   *         ************         *
	5'h11: rom_data2_1234 =  32'b00000000_00000000_00000010_00000001;	//   *                     *        *
	5'h12: rom_data2_1234 =  32'b00000000_00000000_00000011_00000001;	//   *                     **       *
	5'h13: rom_data2_1234 =  32'b00000000_00000000_00000011_00000001;	//   *                     **       *
	5'h14: rom_data2_1234 =  32'b00000000_00000000_00000011_00000001;	//   *                     **       *
	5'h15: rom_data2_1234 =  32'b00000000_00000000_00000011_00000001;	//   *                     **       *
	5'h16: rom_data2_1234 =  32'b00000000_00000000_00000011_00000001;	//   *                     **       *
	5'h17: rom_data2_1234 =  32'b00000000_00000000_00000011_00000001;	//   *                     **       *
	5'h18: rom_data2_1234 =  32'b00000000_00000000_00000011_00000001;	//   *                     **       *
	5'h19: rom_data2_1234 =  32'b00000000_00000000_00000011_00000001;	//   *                     **       *
	5'h1A: rom_data2_1234 =  32'b00000000_00000000_00000010_00000001;	//   *                     *        *
	5'h1B: rom_data2_1234 =  32'b00000000_00111111_11111100_00000001;	//   *         ************         *
	5'h1C: rom_data2_1234 =  32'b00000000_00011111_11111000_00000001;	//   *          **********          *
	5'h1D: rom_data2_1234 =  32'b00000000_00000000_00000000_00000001; 	//   *				    *
	5'h1E: rom_data2_1234 =  32'b00000000_00000000_00000000_00000001; 	//   *				    *
	5'h1F: rom_data2_1234 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr2_1234 = pix_y[4:0] - NUM_y_t_1234[4:0];
assign rom_col2_1234 = pix_x[4:0] - NUM_x_l_1234[4:0];

//------------------------------------//
// Number 3
wire [4:0] rom_addr3_1234, rom_col3_1234;
reg [31:0] rom_data3_1234;

// number image ROM
always @*
case (rom_addr3_1234)
	5'h0: rom_data3_1234 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data3_1234 =   32'b00000000_00000000_00000000_00000001;	//   *                              *
	5'h2: rom_data3_1234 =   32'b00000000_00000000_00000000_00000001;	//   *                              *
	5'h3: rom_data3_1234 =   32'b00000000_00011111_11111000_00000001;	//   *          **********          *
	5'h4: rom_data3_1234 =   32'b00000000_00111111_11111100_00000001;	//   *         ************         *
	5'h5: rom_data3_1234 =   32'b00000000_01000000_00000010_00000001;	//   *        *            *        *
	5'h6: rom_data3_1234 =   32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h7: rom_data3_1234 =   32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h8: rom_data3_1234 =   32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h9: rom_data3_1234 =   32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'hA: rom_data3_1234 =   32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'hB: rom_data3_1234 =   32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'hC: rom_data3_1234 =   32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'hD: rom_data3_1234 =   32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'hE: rom_data3_1234 =   32'b00000000_01000000_00000000_00000001;	//   *        *                     *
	5'hF: rom_data3_1234 =   32'b00000000_00111111_11111100_00000001;	//   *         ************         *
	5'h10: rom_data3_1234 =  32'b00000000_00111111_11111100_00000001; 	//   *         ************         *
	5'h11: rom_data3_1234 =  32'b00000000_01000000_00000000_00000001;	//   *        *                     *
	5'h12: rom_data3_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h13: rom_data3_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h14: rom_data3_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h15: rom_data3_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h16: rom_data3_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h17: rom_data3_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h18: rom_data3_1234 =  32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h19: rom_data3_1234 =  32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h1A: rom_data3_1234 =  32'b00000000_01000000_00000010_00000001;	//   *        *            *        *
	5'h1B: rom_data3_1234 =  32'b00000000_00111111_11111100_00000001;	//   *         ************         *
	5'h1C: rom_data3_1234 =  32'b00000000_00011111_11111000_00000001;	//   *          **********          *
	5'h1D: rom_data3_1234 =  32'b00000000_00000000_00000000_00000001; 	//   *				    *
	5'h1E: rom_data3_1234 =  32'b00000000_00000000_00000000_00000001; 	//   *				    *
	5'h1F: rom_data3_1234 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr3_1234 = pix_y[4:0] - NUM_y_t_1234[4:0];
assign rom_col3_1234 = pix_x[4:0] - NUM_x_l_1234[4:0];

//------------------------------------//
// Number 4
wire [4:0] rom_addr4_1234, rom_col4_1234;
reg [31:0] rom_data4_1234;

// number image ROM
always @*
case (rom_addr4_1234)
	5'h0: rom_data4_1234 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data4_1234 =   32'b00000000_00000000_00000000_00000001;	//   *                              *
	5'h2: rom_data4_1234 =   32'b00000000_00000000_00000000_00000001;	//   *                              *
	5'h3: rom_data4_1234 =   32'b00000000_00000000_00000000_00000001;	//   *                              *
	5'h4: rom_data4_1234 =   32'b00000000_00000000_00000000_00000001;	//   *                              *
	5'h5: rom_data4_1234 =   32'b00000000_01000000_00000010_00000001;	//   *        *            *        *
	5'h6: rom_data4_1234 =   32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h7: rom_data4_1234 =   32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h8: rom_data4_1234 =   32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h9: rom_data4_1234 =   32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'hA: rom_data4_1234 =   32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'hB: rom_data4_1234 =   32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'hC: rom_data4_1234 =   32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'hD: rom_data4_1234 =   32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'hE: rom_data4_1234 =   32'b00000000_01000000_00000010_00000001;	//   *        *            *        *
	5'hF: rom_data4_1234 =   32'b00000000_00111111_11111100_00000001;	//   *         ************         *
	5'h10: rom_data4_1234 =  32'b00000000_00111111_11111100_00000001; 	//   *         ************         *
	5'h11: rom_data4_1234 =  32'b00000000_01000000_00000000_00000001;	//   *        *                     *
	5'h12: rom_data4_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h13: rom_data4_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h14: rom_data4_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h15: rom_data4_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h16: rom_data4_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h17: rom_data4_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h18: rom_data4_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h19: rom_data4_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h1A: rom_data4_1234 =  32'b00000000_01000000_00000000_00000001;	//   *        *                     *
	5'h1B: rom_data4_1234 =  32'b00000000_00000000_00000000_00000001; 	//   *				    *
	5'h1C: rom_data4_1234 =  32'b00000000_00000000_00000000_00000001; 	//   *				    *
	5'h1D: rom_data4_1234 =  32'b00000000_00000000_00000000_00000001; 	//   *				    *
	5'h1E: rom_data4_1234 =  32'b00000000_00000000_00000000_00000001; 	//   *				    *
	5'h1F: rom_data4_1234 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr4_1234 = pix_y[4:0] - NUM_y_t_1234[4:0];
assign rom_col4_1234 = pix_x[4:0] - NUM_x_l_1234[4:0];

//------------------------------------//
// Number 5
wire [4:0] rom_addr5_1234, rom_col5_1234;
reg [31:0] rom_data5_1234;

// number image ROM
always @*
case (rom_addr5_1234)
	5'h0: rom_data5_1234 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data5_1234 =   32'b00000000_00000000_00000000_00000001;	//   *                              *
	5'h2: rom_data5_1234 =   32'b00000000_00000000_00000000_00000001;	//   *                              *
	5'h3: rom_data5_1234 =   32'b00000000_00011111_11111000_00000001;	//   *          **********          *
	5'h4: rom_data5_1234 =   32'b00000000_00111111_11111100_00000001;	//   *         ************         *
	5'h5: rom_data5_1234 =   32'b00000000_00000000_00000010_00000001;	//   *                     *        *
	5'h6: rom_data5_1234 =   32'b00000000_00000000_00000011_00000001;	//   *                     **       *
	5'h7: rom_data5_1234 =   32'b00000000_00000000_00000011_00000001;	//   *                     **       *
	5'h8: rom_data5_1234 =   32'b00000000_00000000_00000011_00000001;	//   *                     **       *
	5'h9: rom_data5_1234 =   32'b00000000_00000000_00000011_00000001;	//   *                     **       *
	5'hA: rom_data5_1234 =   32'b00000000_00000000_00000011_00000001;	//   *                     **       *
	5'hB: rom_data5_1234 =   32'b00000000_00000000_00000011_00000001;	//   *                     **       *
	5'hC: rom_data5_1234 =   32'b00000000_00000000_00000011_00000001;	//   *                     **       *
	5'hD: rom_data5_1234 =   32'b00000000_00000000_00000011_00000001;	//   *                     **       *
	5'hE: rom_data5_1234 =   32'b00000000_00000000_00000010_00000001;	//   *                     *        *
	5'hF: rom_data5_1234 =   32'b00000000_00111111_11111100_00000001;	//   *         ************         *
	5'h10: rom_data5_1234 =  32'b00000000_00111111_11111100_00000001; 	//   *         ************         *
	5'h11: rom_data5_1234 =  32'b00000000_01000000_00000000_00000001;	//   *        *                     *
	5'h12: rom_data5_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h13: rom_data5_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h14: rom_data5_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h15: rom_data5_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h16: rom_data5_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h17: rom_data5_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h18: rom_data5_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h19: rom_data5_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h1A: rom_data5_1234 =  32'b00000000_01000000_00000000_00000001;	//   *        *                     *
	5'h1B: rom_data5_1234 =  32'b00000000_00111111_11111100_00000001;	//   *         ************         *
	5'h1C: rom_data5_1234 =  32'b00000000_00011111_11111000_00000001;	//   *          **********          *
	5'h1D: rom_data5_1234 =  32'b00000000_00000000_00000000_00000001; 	//   *				    *
	5'h1E: rom_data5_1234 =  32'b00000000_00000000_00000000_00000001; 	//   *				    *
	5'h1F: rom_data5_1234 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr5_1234 = pix_y[4:0] - NUM_y_t_1234[4:0];
assign rom_col5_1234 = pix_x[4:0] - NUM_x_l_1234[4:0];

//------------------------------------//
// Number 6
wire [4:0] rom_addr6_1234, rom_col6_1234;
reg [31:0] rom_data6_1234;

// number image ROM
always @*
case (rom_addr6_1234)
	5'h0: rom_data6_1234 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data6_1234 =   32'b00000000_00000000_00000000_00000001;	//   *                              *
	5'h2: rom_data6_1234 =   32'b00000000_00000000_00000000_00000001;	//   *                              *
	5'h3: rom_data6_1234 =   32'b00000000_00011111_11111000_00000001;	//   *          **********          *
	5'h4: rom_data6_1234 =   32'b00000000_00111111_11111100_00000001;	//   *         ************         *
	5'h5: rom_data6_1234 =   32'b00000000_00000000_00000010_00000001;	//   *                     *        *
	5'h6: rom_data6_1234 =   32'b00000000_00000000_00000011_00000001;	//   *                     **       *
	5'h7: rom_data6_1234 =   32'b00000000_00000000_00000011_00000001;	//   *                     **       *
	5'h8: rom_data6_1234 =   32'b00000000_00000000_00000011_00000001;	//   *                     **       *
	5'h9: rom_data6_1234 =   32'b00000000_00000000_00000011_00000001;	//   *                     **       *
	5'hA: rom_data6_1234 =   32'b00000000_00000000_00000011_00000001;	//   *                     **       *
	5'hB: rom_data6_1234 =   32'b00000000_00000000_00000011_00000001;	//   *                     **       *
	5'hC: rom_data6_1234 =   32'b00000000_00000000_00000011_00000001;	//   *                     **       *
	5'hD: rom_data6_1234 =   32'b00000000_00000000_00000011_00000001;	//   *                     **       *
	5'hE: rom_data6_1234 =   32'b00000000_00000000_00000010_00000001;	//   *                     *        *
	5'hF: rom_data6_1234 =   32'b00000000_00111111_11111100_00000001;	//   *         ************         *
	5'h10: rom_data6_1234 =  32'b00000000_00111111_11111100_00000001; 	//   *         ************         *
	5'h11: rom_data6_1234 =  32'b00000000_01000000_00000010_00000001;	//   *        *            *        *
	5'h12: rom_data6_1234 =  32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h13: rom_data6_1234 =  32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h14: rom_data6_1234 =  32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h15: rom_data6_1234 =  32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h16: rom_data6_1234 =  32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h17: rom_data6_1234 =  32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h18: rom_data6_1234 =  32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h19: rom_data6_1234 =  32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h1A: rom_data6_1234 =  32'b00000000_01000000_00000010_00000001;	//   *        *            *        *
	5'h1B: rom_data6_1234 =  32'b00000000_00111111_11111100_00000001;	//   *         ************         *
	5'h1C: rom_data6_1234 =  32'b00000000_00011111_11111000_00000001;	//   *          **********          *
	5'h1D: rom_data6_1234 =  32'b00000000_00000000_00000000_00000001; 	//   *				    *
	5'h1E: rom_data6_1234 =  32'b00000000_00000000_00000000_00000001; 	//   *				    *
	5'h1F: rom_data6_1234 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr6_1234 = pix_y[4:0] - NUM_y_t_1234[4:0];
assign rom_col6_1234 = pix_x[4:0] - NUM_x_l_1234[4:0];

//------------------------------------//
// Number 7
wire [4:0] rom_addr7_1234, rom_col7_1234;
reg [31:0] rom_data7_1234;

// number image ROM
always @*
case (rom_addr7_1234)
	5'h0: rom_data7_1234 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data7_1234 =   32'b00000000_00000000_00000000_00000001;	//   *                              *
	5'h2: rom_data7_1234 =   32'b00000000_00000000_00000000_00000001;	//   *                              *
	5'h3: rom_data7_1234 =   32'b00000000_00011111_11111000_00000001;	//   *          **********          *
	5'h4: rom_data7_1234 =   32'b00000000_00111111_11111100_00000001;	//   *         ************         *
	5'h5: rom_data7_1234 =   32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h6: rom_data7_1234 =   32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h7: rom_data7_1234 =   32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h8: rom_data7_1234 =   32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h9: rom_data7_1234 =   32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'hA: rom_data7_1234 =   32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'hB: rom_data7_1234 =   32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'hC: rom_data7_1234 =   32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'hD: rom_data7_1234 =   32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'hE: rom_data7_1234 =   32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'hF: rom_data7_1234 =   32'b00000000_01000000_00000000_00000001;	//   *        *                     *
	5'h10: rom_data7_1234 =  32'b00000000_01000000_00000000_00000001;	//   *        *                     *
	5'h11: rom_data7_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h12: rom_data7_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h13: rom_data7_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h14: rom_data7_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h15: rom_data7_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h16: rom_data7_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h17: rom_data7_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h18: rom_data7_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h19: rom_data7_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h1A: rom_data7_1234 =  32'b00000000_01000000_00000000_00000001;	//   *        *                     *
	5'h1B: rom_data7_1234 =  32'b00000000_00000000_00000000_00000001; 	//   *				    *
	5'h1C: rom_data7_1234 =  32'b00000000_00000000_00000000_00000001; 	//   *				    *
	5'h1D: rom_data7_1234 =  32'b00000000_00000000_00000000_00000001; 	//   *				    *
	5'h1E: rom_data7_1234 =  32'b00000000_00000000_00000000_00000001; 	//   *				    *
	5'h1F: rom_data7_1234 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr7_1234 = pix_y[4:0] - NUM_y_t_1234[4:0];
assign rom_col7_1234 = pix_x[4:0] - NUM_x_l_1234[4:0];

//------------------------------------//
// Number 8
wire [4:0] rom_addr8_1234, rom_col8_1234;
reg [31:0] rom_data8_1234;

// number image ROM
always @*
case (rom_addr8_1234)
	5'h0: rom_data8_1234 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data8_1234 =   32'b00000000_00000000_00000000_00000001;	//   *                              *
	5'h2: rom_data8_1234 =   32'b00000000_00000000_00000000_00000001;	//   *                              *
	5'h3: rom_data8_1234 =   32'b00000000_00011111_11111000_00000001;	//   *          **********          *
	5'h4: rom_data8_1234 =   32'b00000000_00111111_11111100_00000001;	//   *         ************         *
	5'h5: rom_data8_1234 =   32'b00000000_01000000_00000010_00000001;	//   *        *            *        *
	5'h6: rom_data8_1234 =   32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h7: rom_data8_1234 =   32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h8: rom_data8_1234 =   32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h9: rom_data8_1234 =   32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'hA: rom_data8_1234 =   32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'hB: rom_data8_1234 =   32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'hC: rom_data8_1234 =   32'b00000000_11000000_00000011_00000000;	//   *       **            **       *
	5'hD: rom_data8_1234 =   32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'hE: rom_data8_1234 =   32'b00000000_01000000_00000010_00000001;	//   *        *            *        *
	5'hF: rom_data8_1234 =   32'b00000000_00111111_11111100_00000001;	//   *         ************         *
	5'h10: rom_data8_1234 =  32'b00000000_00111111_11111100_00000001; 	//   *         ************         *
	5'h11: rom_data8_1234 =  32'b00000000_01000000_00000010_00000001;	//   *        *            *        *
	5'h12: rom_data8_1234 =  32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h13: rom_data8_1234 =  32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h14: rom_data8_1234 =  32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h15: rom_data8_1234 =  32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h16: rom_data8_1234 =  32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h17: rom_data8_1234 =  32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h18: rom_data8_1234 =  32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h19: rom_data8_1234 =  32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h1A: rom_data8_1234 =  32'b00000000_01000000_00000010_00000001;	//   *        *            *        *
	5'h1B: rom_data8_1234 =  32'b00000000_00111111_11111100_00000001;	//   *         ************         *
	5'h1C: rom_data8_1234 =  32'b00000000_00011111_11111000_00000001;	//   *          **********          *
	5'h1D: rom_data8_1234 =  32'b00000000_00000000_00000000_00000001; 	//   *				    *
	5'h1E: rom_data8_1234 =  32'b00000000_00000000_00000000_00000001; 	//   *				    *
	5'h1F: rom_data8_1234 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr8_1234 = pix_y[4:0] - NUM_y_t_1234[4:0];
assign rom_col8_1234 = pix_x[4:0] - NUM_x_l_1234[4:0];

//------------------------------------//
// Number 9
wire [4:0] rom_addr9_1234, rom_col9_1234;
reg [31:0] rom_data9_1234;

// number image ROM
always @*
case (rom_addr9_1234)
	5'h0: rom_data9_1234 =   32'b11111111_11111111_11111111_11111111;	//   ********************************
	5'h1: rom_data9_1234 =   32'b00000000_00000000_00000000_00000001;	//   *                              *
	5'h2: rom_data9_1234 =   32'b00000000_00000000_00000000_00000001;	//   *                              *
	5'h3: rom_data9_1234 =   32'b00000000_00011111_11111000_00000001;	//   *          **********          *
	5'h4: rom_data9_1234 =   32'b00000000_00111111_11111100_00000001;	//   *         ************         *
	5'h5: rom_data9_1234 =   32'b00000000_01000000_00000010_00000001;	//   *        *            *        *
	5'h6: rom_data9_1234 =   32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h7: rom_data9_1234 =   32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h8: rom_data9_1234 =   32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'h9: rom_data9_1234 =   32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'hA: rom_data9_1234 =   32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'hB: rom_data9_1234 =   32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'hC: rom_data9_1234 =   32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'hD: rom_data9_1234 =   32'b00000000_11000000_00000011_00000001;	//   *       **            **       *
	5'hE: rom_data9_1234 =   32'b00000000_01000000_00000010_00000001;	//   *        *            *        *
	5'hF: rom_data9_1234 =   32'b00000000_00111111_11111100_00000001;	//   *         ************         *
	5'h10: rom_data9_1234 =  32'b00000000_00111111_11111100_00000001; 	//   *         ************         *
	5'h11: rom_data9_1234 =  32'b00000000_01000000_00000000_00000001;	//   *        *                     *
	5'h12: rom_data9_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h13: rom_data9_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h14: rom_data9_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h15: rom_data9_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h16: rom_data9_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h17: rom_data9_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h18: rom_data9_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h19: rom_data9_1234 =  32'b00000000_11000000_00000000_00000001;	//   *       **                     *
	5'h1A: rom_data9_1234 =  32'b00000000_01000000_00000000_00000001;	//   *        *                     *
	5'h1B: rom_data9_1234 =  32'b00000000_00000000_00000000_00000001; 	//   *				    *
	5'h1C: rom_data9_1234 =  32'b00000000_00000000_00000000_00000001; 	//   *				    *
	5'h1D: rom_data9_1234 =  32'b00000000_00000000_00000000_00000001; 	//   *				    *
	5'h1E: rom_data9_1234 =  32'b00000000_00000000_00000000_00000001; 	//   *				    *
	5'h1F: rom_data9_1234 =  32'b11111111_11111111_11111111_11111111;	//   ********************************
endcase

// Map current pixel location to ROM addr/col
assign rom_addr9_1234 = pix_y[4:0] - NUM_y_t_1234[4:0];
assign rom_col9_1234 = pix_x[4:0] - NUM_x_l_1234[4:0];

always @(posedge clk) begin
	if (score[15:12] == 0)
	    rom_bit_1234 = rom_data0_1234[rom_col0_1234];
	else if (score[15:12] == 1)
	    rom_bit_1234 = rom_data1_1234[rom_col1_1234];
	else if (score[15:12] == 2)
	    rom_bit_1234 = rom_data2_1234[rom_col2_1234];
	else if (score[15:12] == 3)
	    rom_bit_1234 = rom_data3_1234[rom_col3_1234];
	else if (score[15:12] == 4)
	    rom_bit_1234 = rom_data4_1234[rom_col4_1234];
	else if (score[15:12] == 5)
	    rom_bit_1234 = rom_data5_1234[rom_col5_1234];
	else if (score[15:12] == 6)
	    rom_bit_1234 = rom_data6_1234[rom_col6_1234];
	else if (score[15:12] == 7)
	    rom_bit_1234 = rom_data7_1234[rom_col7_1234];
	else if (score[15:12] == 8)
	    rom_bit_1234 = rom_data8_1234[rom_col8_1234];
	else if (score[15:12] == 9)
	    rom_bit_1234 = rom_data9_1234[rom_col9_1234];
end


// Pixel within a block
assign NUM_one =  ((NUM_x_l_1 <= pix_x) && (pix_x <= NUM_x_r_1) && (NUM_y_t_1 <= pix_y) && (pix_y <= NUM_y_b_1));  
assign NUM_two = ((NUM_x_l_12 <= pix_x) && (pix_x <= NUM_x_r_12) && (NUM_y_t_12 <= pix_y) && (pix_y <= NUM_y_b_12)); 
assign NUM_three = ((NUM_x_l_123 <= pix_x) && (pix_x <= NUM_x_r_123) && (NUM_y_t_123 <= pix_y) && (pix_y <= NUM_y_b_123));
assign NUM_four = ((NUM_x_l_1234 <= pix_x) && (pix_x <= NUM_x_r_1234) && (NUM_y_t_1234 <= pix_y) && (pix_y <= NUM_y_b_1234));

// Pixel within number
assign score_ON_R = NUM_one && rom_bit_1;
assign score_ON_RM = NUM_two && rom_bit_12;
assign score_ON_LM = NUM_three && rom_bit_123;
assign score_ON_L = NUM_four && rom_bit_1234;

endmodule
